module rotate_left(input wire [31:0] a, b, output wire [31:0] result);
begin
	wire [4:0] bits;
	
end